library verilog;
use verilog.vl_types.all;
entity lab7 is
    port(
        S0              : out    vl_logic;
        C0              : in     vl_logic;
        x0              : in     vl_logic;
        y0              : in     vl_logic;
        S1              : out    vl_logic;
        x1              : in     vl_logic;
        y1              : in     vl_logic;
        S2              : out    vl_logic;
        x2              : in     vl_logic;
        y2              : in     vl_logic;
        S3              : out    vl_logic;
        x3              : in     vl_logic;
        y3              : in     vl_logic;
        C3              : out    vl_logic;
        S4              : out    vl_logic
    );
end lab7;
