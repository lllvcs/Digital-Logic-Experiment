library verilog;
use verilog.vl_types.all;
entity lab8 is
    port(
        Q3              : out    vl_logic;
        CLK             : in     vl_logic;
        D               : in     vl_logic;
        Q4              : out    vl_logic;
        K               : in     vl_logic;
        J               : in     vl_logic;
        Q5              : out    vl_logic;
        T               : in     vl_logic;
        Q1              : out    vl_logic;
        R               : in     vl_logic;
        S               : in     vl_logic;
        Q2              : out    vl_logic;
        NR              : in     vl_logic;
        NS              : in     vl_logic;
        NQ1             : out    vl_logic;
        NQ2             : out    vl_logic
    );
end lab8;
