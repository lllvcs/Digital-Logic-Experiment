library verilog;
use verilog.vl_types.all;
entity lab7_vlg_vec_tst is
end lab7_vlg_vec_tst;
