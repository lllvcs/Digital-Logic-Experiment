library verilog;
use verilog.vl_types.all;
entity lab8_vlg_vec_tst is
end lab8_vlg_vec_tst;
