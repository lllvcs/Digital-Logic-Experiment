library verilog;
use verilog.vl_types.all;
entity lab9_vlg_vec_tst is
end lab9_vlg_vec_tst;
