library verilog;
use verilog.vl_types.all;
entity lab9_vlg_check_tst is
    port(
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        c1              : in     vl_logic;
        c2              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        e1              : in     vl_logic;
        e2              : in     vl_logic;
        f1              : in     vl_logic;
        f2              : in     vl_logic;
        g1              : in     vl_logic;
        g2              : in     vl_logic;
        Q11             : in     vl_logic;
        Q12             : in     vl_logic;
        Q13             : in     vl_logic;
        Q14             : in     vl_logic;
        Q21             : in     vl_logic;
        Q22             : in     vl_logic;
        Q23             : in     vl_logic;
        Q24             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab9_vlg_check_tst;
