library verilog;
use verilog.vl_types.all;
entity lab8_vlg_check_tst is
    port(
        NQ1             : in     vl_logic;
        NQ2             : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        Q3              : in     vl_logic;
        Q4              : in     vl_logic;
        Q5              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab8_vlg_check_tst;
