library verilog;
use verilog.vl_types.all;
entity lab11 is
    port(
        a1              : out    vl_logic;
        pin7            : in     vl_logic;
        a2              : out    vl_logic;
        a3              : out    vl_logic;
        a4              : out    vl_logic;
        a5              : out    vl_logic;
        a6              : out    vl_logic;
        a               : out    vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic
    );
end lab11;
