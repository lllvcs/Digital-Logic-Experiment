library verilog;
use verilog.vl_types.all;
entity lab6_3_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Ci_1            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab6_3_vlg_sample_tst;
