library verilog;
use verilog.vl_types.all;
entity lab11_vlg_vec_tst is
end lab11_vlg_vec_tst;
