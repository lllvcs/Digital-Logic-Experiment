library verilog;
use verilog.vl_types.all;
entity ex2_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ex2_vlg_check_tst;
