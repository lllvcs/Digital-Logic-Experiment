library verilog;
use verilog.vl_types.all;
entity lab11_vlg_sample_tst is
    port(
        pin7            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab11_vlg_sample_tst;
