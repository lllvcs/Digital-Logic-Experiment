library verilog;
use verilog.vl_types.all;
entity lab6_3_vlg_check_tst is
    port(
        Ci              : in     vl_logic;
        Si              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab6_3_vlg_check_tst;
