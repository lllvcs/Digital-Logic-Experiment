library verilog;
use verilog.vl_types.all;
entity lab6_3 is
    port(
        Si              : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        Ci_1            : in     vl_logic;
        Ci              : out    vl_logic
    );
end lab6_3;
