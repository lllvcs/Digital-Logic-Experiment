library verilog;
use verilog.vl_types.all;
entity lab10_vlg_vec_tst is
end lab10_vlg_vec_tst;
