library verilog;
use verilog.vl_types.all;
entity lab9 is
    port(
        Q11             : out    vl_logic;
        CLK             : in     vl_logic;
        Q12             : out    vl_logic;
        Q13             : out    vl_logic;
        Q14             : out    vl_logic;
        a1              : out    vl_logic;
        b1              : out    vl_logic;
        c1              : out    vl_logic;
        d1              : out    vl_logic;
        e1              : out    vl_logic;
        f1              : out    vl_logic;
        g1              : out    vl_logic;
        a2              : out    vl_logic;
        b2              : out    vl_logic;
        c2              : out    vl_logic;
        d2              : out    vl_logic;
        e2              : out    vl_logic;
        f2              : out    vl_logic;
        g2              : out    vl_logic;
        Q24             : out    vl_logic;
        Q23             : out    vl_logic;
        Q21             : out    vl_logic;
        Q22             : out    vl_logic
    );
end lab9;
