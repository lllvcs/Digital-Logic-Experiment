library verilog;
use verilog.vl_types.all;
entity extra_vlg_vec_tst is
end extra_vlg_vec_tst;
